`default_nettype none

module abstractChipInterface();
endmodule:abstractChipInterface
